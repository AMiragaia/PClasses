library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity fsm is
		port(reset 		 : in std_logic;
			  start      : in std_logic;
			  clk   		 : in std_logic;
			  filter_on  : in std_logic;
			  rst_ram	 :	in std_logic;
			  algarismo1 : out std_logic_vector(6 downto 0);
			  algarismo2 : out std_logic_vector(6 downto 0);
			  algarismo3 : out std_logic_vector(6 downto 0);
			  algarismo4 : out std_logic_vector(6 downto 0);
			  algarismo5 : out std_logic_vector(6 downto 0);
			  algarismo6 : out std_logic_vector(6 downto 0);
			  algarismo7 : out std_logic_vector(6 downto 0);
			  algarismo8 : out std_logic_vector(6 downto 0));

architecture Behavioral of fsm is
	
			  
			  
			  