library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity NoisyTriangSignal_ROM_256x8 is
   port(address : in  std_logic_vector(7 downto 0);
        dataOut : out std_logic_vector(7 downto 0));
end NoisyTriangSignal_ROM_256x8;

architecture Behavioral of NoisyTriangSignal_ROM_256x8 is
   subtype TDataWord is std_logic_vector(7 downto 0);
   type TROM is array (0 to 255) of TDataWord;
	-- Input Signal ROM
   constant c_memory: TROM := (
	"10101001",
	"10101101",
	"10010010",
	"10101001",
	"10100100",
	"10101011",
	"11000100",
	"10101111",
	"10101001",
	"10111110",
	"10111111",
	"10111111",
	"11001111",
	"11001111",
	"11010000",
	"11001101",
	"11010111",
	"11010100",
	"11011011",
	"11100010",
	"11100011",
	"11011101",
	"11100001",
	"11100000",
	"11110110",
	"11110000",
	"11101101",
	"11111101",
	"11110101",
	"00000001",
	"00001111",
	"00001100",
	"00000101",
	"00001001",
	"00011111",
	"00001110",
	"00010110",
	"00011010",
	"00100010",
	"00011111",
	"00100100",
	"00100110",
	"01000000",
	"00110010",
	"00100100",
	"00100100",
	"00100100",
	"01001000",
	"00110010",
	"01000110",
	"01000101",
	"00110101",
	"01011010",
	"01001111",
	"01011110",
	"01010011",
	"01010101",
	"01001101",
	"01011010",
	"01011110",
	"01010001",
	"01011101",
	"01011011",
	"01001111",
	"01010111",
	"01000100",
	"01000111",
	"01001011",
	"01000001",
	"01000111",
	"00111101",
	"00110100",
	"01000011",
	"00111100",
	"00111001",
	"00110111",
	"00110110",
	"00110011",
	"00100111",
	"00011111",
	"00011111",
	"00101001",
	"00001110",
	"00010001",
	"00011101",
	"00011000",
	"00001000",
	"00001000",
	"00000101",
	"00000001",
	"11101001",
	"11111001",
	"11111101",
	"00001110",
	"11100101",
	"11101010",
	"11101001",
	"11100001",
	"11100000",
	"11010001",
	"11011111",
	"11011000",
	"11011111",
	"11010111",
	"11011101",
	"11100000",
	"11001110",
	"10111110",
	"11001001",
	"11010001",
	"10111111",
	"11000001",
	"10110000",
	"11000101",
	"10110111",
	"10101100",
	"10011101",
	"10100011",
	"10011101",
	"10011110",
	"10100011",
	"10101011",
	"10101000",
	"10101010",
	"10110000",
	"11001001",
	"10110110",
	"10111000",
	"11001001",
	"10111110",
	"10111010",
	"11001100",
	"11000011",
	"11001100",
	"11010101",
	"11011000",
	"11000100",
	"11000000",
	"11010011",
	"11101101",
	"11100010",
	"11100010",
	"11100101",
	"11110100",
	"11110000",
	"11110101",
	"11011111",
	"11110101",
	"11111010",
	"11110101",
	"00000000",
	"11111101",
	"00001111",
	"00000100",
	"00011001",
	"00010000",
	"00011100",
	"00101100",
	"00011010",
	"00101011",
	"00010110",
	"00110101",
	"00011011",
	"00101001",
	"00101010",
	"00100101",
	"00100111",
	"00111101",
	"00101100",
	"00110000",
	"01001011",
	"01000011",
	"01001010",
	"01000001",
	"01001011",
	"01010011",
	"01010101",
	"01101000",
	"01010100",
	"01011011",
	"01101000",
	"01100110",
	"01000111",
	"01010011",
	"01001101",
	"01010000",
	"01010010",
	"01001110",
	"01010001",
	"01000111",
	"01000011",
	"01000110",
	"00111110",
	"00101010",
	"00110100",
	"00100000",
	"00110111",
	"00010101",
	"00100001",
	"00100100",
	"00100000",
	"00101111",
	"00011010",
	"00010001",
	"00011001",
	"00000100",
	"00010010",
	"00001100",
	"00000011",
	"11111101",
	"11110101",
	"11101011",
	"11110110",
	"11111110",
	"11101100",
	"11111111",
	"11100100",
	"11111110",
	"11100000",
	"11100100",
	"11101110",
	"11101001",
	"11010010",
	"11011101",
	"11001001",
	"11000000",
	"11010011",
	"10111001",
	"10110010",
	"11000011",
	"11001101",
	"11001000",
	"10101011",
	"10110111",
	"10111011",
	"10111001",
	"10111100",
	"10111001",
	"10101111",
	"10010110",
	"10100000",
	"10010110",
	"10110010",
	"10111010",
	"10011010",
	"10111000",
	"10110000",
	"10110010",
	"10110001",
	"11001001",
	"11000100",
	"11000010",
	"11001010",
	"11010011",
	"11000100",
	"11001000");

begin
   dataOut <= c_memory(to_integer(unsigned(address)));
end Behavioral;




