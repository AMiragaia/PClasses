library ieee;
use ieee.std_logic_1164.all;

entity dec4_16 is
	port(inputs : in std_logic_vector(3 downto 0);
		  outputs : out std_logic_vector(15 downto 0));
end dec4_16;


--decoder feito para valor decimal aparecer na led respetiva
architecture behavioral of dec4_16 is
begin
	process(inputs)
	begin
		 case inputs is
		 when "0000" =>
		 outputs <= "0000000000000001";
		 when "0001" =>
		 outputs <= "0000000000000010";
		 when "0010" =>
		 outputs <= "0000000000000100";
		 when "0011" =>
		 outputs <= "0000000000001000";
		 when "0100" =>
		 outputs <= "0000000000010000";
		 when "0101" =>
		 outputs <= "0000000000100000";
		 when "0110" =>
		 outputs <= "0000000001000000";
		 when "0111" =>
		 outputs <= "0000000010000000";
		 when "1000" =>
		 outputs <= "0000000100000000";
		 when "1001" =>
		 outputs <= "0000001000000000";
		 when "1010" =>
		 outputs <= "0000010000000000";
		 when "1011" =>
		 outputs <= "0000100000000000";
		 when "1100" =>
		 outputs <= "0001000000000000";
		 when "1101" =>
		 outputs <= "0010000000000000";
		 when "1110" =>
		 outputs <= "0100000000000000";
		 when "1111" =>
		 outputs <= "1000000000000000";
		 when others =>
		 outputs <= "0000000000000000";
		 end case;
		
	end process;
end Behavioral;
